  UILANG="Svenska"  
  label="ID (uid/gid)"  
  label_homeDir="Hemkatalog"  
  label_loginShell="Inloggningsskal"  
  label_realName="Riktigt namn"  
  label_room="Rum"  
  label_workPhone="Arbetstelefon"  
  label_phone="Hemtelefon"  
  label_comment="Kommentar"
  
  field_descriptions[1]="Användarnamn;Inloggningsnamn för användaren;namn"
  field_descriptions[2]="Lösenord;Platshållare för krypterat lösenord (vanligtvis 'x')"
  field_descriptions[3]="UID;Användar-ID-nummer"
  field_descriptions[4]="GID;Primärt grupp-ID-nummer"
  field_descriptions[5]="GECOS;Användarinformation (fullständigt namn, kontaktuppgifter)"
  field_descriptions[6]="Hemkatalog;Sökväg till användarens hemkatalog;katalog"
  field_descriptions[7]="Inloggningsskal;Sökväg till användarens standardskal;skal"
  
ERROR="FEL"
ERR_INCORRECT_FIELD="Fel namn eller nummer för fält angivet"
INFO_CORRECT_FIELDS="Vänligen använd ett giltigt fältnamn eller fältnummer!"
AVAILABLE_FIELD_NAMES="Tillgängliga fältnamn"
AVAILABLE_FIELD_NUMBERS="Tillgängliga fältnummer"

FIELD="Datfält"
